LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity game_logic is
	generic(
	);
	port(
		
	);
end;

architecture game_logic_bhv of game_logic is
	
begin
	
end;
	
	
