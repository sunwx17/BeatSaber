LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity beatsaber is
	generic(
	);
	port(
	);
end;

architecture main of beatsaber is
	
begin
	
end;
	
	
